module freq_div(clk_in, reset, clk_out);
	parameter exp = 20;   
	input clk_in, reset;
	output clk_out;
	reg[exp-1:0] divider;
	integer i;
	assign clk_out= divider[exp-1];
	always@ (posedge clk_in or posedge reset)	begin
	if(reset)
		for(i=0; i < exp; i=i+1)
			divider[i] = 1'b0;
	else
		divider = divider+ 1'b1;
	end
endmodule 