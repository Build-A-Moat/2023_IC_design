module		map(addr,data);
	input		[5:0]addr;
	output reg 	[7:0]data;
	always@(addr) begin
		case(addr)
			6'd0  :data=8'b0011_1100;
			6'd1  :data=8'b0100_0010;
			6'd2	:data=8'b1010_0101;
			6'd3	:data=8'b1001_1001;
			6'd4	:data=8'b1000_0001;
			6'd5	:data=8'b1010_0101;
			6'd6	:data=8'b0100_0010;
			6'd7	:data=8'b0011_1100;
			
			6'd8  :data=8'b0000_0001;            
			6'd9  :data=8'b0000_0010; 
			6'd10 :data=8'b0000_1100;
			6'd11 :data=8'b0000_0000;
			6'd12 :data=8'b0001_0000;
			6'd13 :data=8'b0010_0000;
			6'd14 :data=8'b0100_0000;
			6'd15 :data=8'b1000_0000;
			
			6'd16 :data=8'b0000_0000;
			6'd17 :data=8'b0000_0000;
			6'd18	:data=8'b0100_0000;
			6'd19	:data=8'b0000_0000;
			6'd20	:data=8'b0011_0000;
			6'd21	:data=8'b0000_1000;
			6'd22	:data=8'b0000_0000;
			6'd23	:data=8'b0000_0000;
			
			6'd24 :data=8'b0000_0100;
			6'd25 :data=8'b0000_1000;
			6'd26	:data=8'b0100_0000;
			6'd27	:data=8'b0000_0000;
			6'd28	:data=8'b0011_0000;
			6'd29	:data=8'b0000_1000;
			6'd30	:data=8'b0000_0000;
			6'd31	:data=8'b0000_0000;
			
			6'd24 :data=8'b0000_0100;
			6'd25 :data=8'b0000_1000;
			6'd26	:data=8'b0100_0000;
			6'd27	:data=8'b0000_0000;
			6'd28	:data=8'b0011_0000;
			6'd29	:data=8'b0000_1000;
			6'd30	:data=8'b0000_0000;
			6'd31	:data=8'b0000_0000;
			
			6'd32 :data=8'b0000_0100;
			6'd33 :data=8'b0001_0000;
			6'd34	:data=8'b0100_0000;
			6'd35	:data=8'b0000_0000;
			6'd36	:data=8'b0011_0000;
			6'd37	:data=8'b0000_1000;
			6'd38	:data=8'b0000_0000;
			6'd39	:data=8'b0000_0000;
			
			6'd40 :data=8'b0000_0100;
			6'd41 :data=8'b0000_1000;
			6'd42	:data=8'b0100_0000;
			6'd43	:data=8'b0000_0000;
			6'd44	:data=8'b0011_0000;
			6'd45	:data=8'b0000_1000;
			6'd46	:data=8'b0000_0000;
			6'd47	:data=8'b0000_0000;
			
			6'd48 :data=8'b0000_0100;
			6'd49 :data=8'b0000_1000;
			6'd50	:data=8'b0100_0000;
			6'd51	:data=8'b0000_0000;
			6'd52	:data=8'b0011_0000;
			6'd53	:data=8'b0000_1000;
			6'd54	:data=8'b0000_0000;
			6'd55	:data=8'b0000_0000;
			
			6'd56 :data=8'b0000_0100;
			6'd57 :data=8'b0000_1000;
			6'd58	:data=8'b0100_0000;
			6'd59 :data=8'b0000_0000;
			6'd60	:data=8'b0000_0000;
			6'd61	:data=8'b0000_0000;
			6'd62	:data=8'b0000_0000;
			6'd63	:data=8'b0000_0000;
			default	:data=8'b0000_0000;
		endcase
	end
endmodule

